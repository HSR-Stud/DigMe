-- Required libraries for ''numeric_std'' implementation
library ieee;
use ieee.numeric_std.all;
use ieee.math_real.all;
-- Required libraries for ''fixed_pkg'' implementation in VHDL 2008
Library ieee;
use ieee.fixed_pkg.all;
use ieee.fixed_float_types.all;
-- Required libraries for ''fixed_pkg'' implementation in older VHDL versions
Library ieee_proposed;
use ieee_proposed.fixed_pkg.all;
use ieee_proposed,fixed_float_types.all;
